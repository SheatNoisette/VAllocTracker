module main

fn main() {
	println('Hello, world!')
	// Print allocations
	custom_alloc_print_stats()
}
